--Modified for the FELIX HTG-710,   Kai CHEN @ bnl 

------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.7
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gth_quad_4p8g_cpll_exdes.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gth_quad_4p8g_cpll_exdes
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity gth_quad_4p8g_cpll_exdes is
generic
(
   
    STABLE_CLOCK_PERIOD                     : integer   := 24

);
port
(
-------------------------------------
---	CLK ---------------------------
-------------------------------------
	 q2_clk0_refclk_in							: in   std_logic; 
    DRP_CLK_IN                            : in   std_logic;
	 
	 --- RX clock, for each channel
	 gt0_rxusrclk_in  : in   std_logic;
	 gt0_rxoutclk_out : out  std_logic;
	 
	 gt1_rxusrclk_in  : in   std_logic;
	 gt1_rxoutclk_out : out  std_logic;
	 
	 gt2_rxusrclk_in  : in   std_logic;
	 gt2_rxoutclk_out : out  std_logic;
	 
	 gt3_rxusrclk_in  : in   std_logic;
	 gt3_rxoutclk_out : out  std_logic;
	 
	 --- TX clock, shared by all channels
	 gt0_txusrclk_in	: in   std_logic;
	 gt0_txoutclk_out : out  std_logic;

-----------------------------------------
---- STATUS signals
-----------------------------------------
	 gt_txresetdone_out   : out  std_logic_vector(3 downto 0); 
    gt_rxresetdone_out   : out  std_logic_vector(3 downto 0);
     
	 gt_txfsmresetdone_out : out  std_logic_vector(3 downto 0);
	 gt_rxfsmresetdone_out : out  std_logic_vector(3 downto 0);
	 
	 gt_cpllfbclklost_out 	: out  std_logic_vector(3 downto 0);
	 gt_cplllock_out 			: out  std_logic_vector(3 downto 0);
	 
	 gt_rxcdrlock_out 		: out  std_logic_vector(3 downto 0);
	 gt_qplllock_out 			: out  std_logic;
---------------------------
---- CTRL signals
---------------------------
	 gt_rxslide_in 			: in   std_logic_vector(3 downto 0);
	 gt_txuserrdy_in       	: in   std_logic_vector(3 downto 0); 
	 gt_rxuserrdy_in       	: in   std_logic_vector(3 downto 0);
	 
----------------------------------------------------------------
----------RESET SIGNALs
----------------------------------------------------------------	 
	 
	 SOFT_RESET_IN 								  : in 	std_logic; 
    GTTX_RESET_IN                           : in   std_logic_vector(3 downto 0);
    GTRX_RESET_IN                           : in   std_logic_vector(3 downto 0);
    CPLL_RESET_IN                           : in   std_logic_vector(3 downto 0);
    QPLL_RESET_IN                           : in   std_logic;
    
     SOFT_TXRST_GT      : in   std_logic_vector(3 downto 0);
       SOFT_RXRST_GT     : in   std_logic_vector(3 downto 0);
       SOFT_TXRST_ALL      : in   std_logic;
       SOFT_RXRST_ALL      : in   std_logic;

-----------------------------------------------------------
----------- Data and TX/RX Ports
-----------------------------------------------------------
	 
	 RX_DATA_gt0_20b : out std_logic_vector(19 downto 0);
	 TX_DATA_gt0_20b : in std_logic_vector(19 downto 0);
	 RX_DATA_gt1_20b : out std_logic_vector(19 downto 0);
	 TX_DATA_gt1_20b : in std_logic_vector(19 downto 0);
	 RX_DATA_gt2_20b : out std_logic_vector(19 downto 0);
	 TX_DATA_gt2_20b : in std_logic_vector(19 downto 0);
	 RX_DATA_gt3_20b : out std_logic_vector(19 downto 0);
	 TX_DATA_gt3_20b : in std_logic_vector(19 downto 0);
	 
    RXN_IN                                  : in   std_logic_vector(3 downto 0);
    RXP_IN                                  : in   std_logic_vector(3 downto 0);
    TXN_OUT                                 : out  std_logic_vector(3 downto 0);
    TXP_OUT                                 : out  std_logic_vector(3 downto 0)
);


end gth_quad_4p8g_cpll_exdes;
    
architecture RTL of gth_quad_4p8g_cpll_exdes is
    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gth_quad_4p8g_cpll_20141208,gtwizard_v2_7,{protocol_file=Start_from_scratch}";

--**************************Component Declarations*****************************

--component gth_quad_4p8g_cpll_init
--generic
--(
--    -- Simulation attributes
--    EXAMPLE_SIM_GTRESET_SPEEDUP    : string    := "FALSE";    -- Set to 1 to speed up sim reset
--    EXAMPLE_SIMULATION             : integer   := 0;          -- Set to 1 for simulation
--    STABLE_CLOCK_PERIOD            : integer   := 6;    --Period of the stable clock driving this state-machine, unit is [ns]
--    EXAMPLE_USE_CHIPSCOPE          : integer   := 0           -- Set to 1 to use Chipscope to drive resets
--);
--port
--(
--    SYSCLK_IN                               : in   std_logic;
--    SOFT_RESET_IN                           : in   std_logic;
--    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
--    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT0_DATA_VALID_IN                       : in   std_logic;
--    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT1_DATA_VALID_IN                       : in   std_logic;
--    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT2_DATA_VALID_IN                       : in   std_logic;
--    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
--    GT3_DATA_VALID_IN                       : in   std_logic;
--
--    --_________________________________________________________________________
--    --_________________________________________________________________________
--    --GT0  (X1Y4)
--    --____________________________CHANNEL PORTS________________________________
--    --------------------------------- CPLL Ports -------------------------------
--    GT0_CPLLFBCLKLOST_OUT                   : out  std_logic;
--    GT0_CPLLLOCK_OUT                        : out  std_logic;
--    GT0_CPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT0_CPLLRESET_IN                        : in   std_logic;
--    -------------------------- Channel - Clocking Ports ------------------------
--    GT0_GTREFCLK0_IN                        : in   std_logic;
--    ---------------------------- Channel - DRP Ports  --------------------------
--    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
--    GT0_DRPCLK_IN                           : in   std_logic;
--    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
--    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
--    GT0_DRPEN_IN                            : in   std_logic;
--    GT0_DRPRDY_OUT                          : out  std_logic;
--    GT0_DRPWE_IN                            : in   std_logic;
--    --------------------- RX Initialization and Reset Ports --------------------
--    GT0_RXUSERRDY_IN                        : in   std_logic;
--    -------------------------- RX Margin Analysis Ports ------------------------
--    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
--    ------------------------- Receive Ports - CDR Ports ------------------------
--    GT0_RXCDRLOCK_OUT                       : out  std_logic;
--    --------------- Receive Ports - Comma Detection and Alignment --------------
--    GT0_RXSLIDE_IN                          : in   std_logic;
--    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--    GT0_RXUSRCLK_IN                         : in   std_logic;
--    GT0_RXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Receive Ports - FPGA RX interface Ports -----------------
--    GT0_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
--    ------------------------ Receive Ports - RX AFE Ports ----------------------
--    GT0_GTHRXN_IN                           : in   std_logic;
--    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--    GT0_RXPHMONITOR_OUT                     : out  std_logic_vector(4 downto 0);
--    GT0_RXPHSLIPMONITOR_OUT                 : out  std_logic_vector(4 downto 0);
--    --------------- Receive Ports - RX Fabric Output Control Ports -------------
--    GT0_RXOUTCLK_OUT                        : out  std_logic;
--    ------------- Receive Ports - RX Initialization and Reset Ports ------------
--    GT0_GTRXRESET_IN                        : in   std_logic;
--    ------------------------ Receive Ports -RX AFE Ports -----------------------
--    GT0_GTHRXP_IN                           : in   std_logic;
--    -------------- Receive Ports -RX Initialization and Reset Ports ------------
--    GT0_RXRESETDONE_OUT                     : out  std_logic;
--    --------------------- TX Initialization and Reset Ports --------------------
--    GT0_GTTXRESET_IN                        : in   std_logic;
--    GT0_TXUSERRDY_IN                        : in   std_logic;
--    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--    GT0_TXUSRCLK_IN                         : in   std_logic;
--    GT0_TXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Transmit Ports - TX Data Path interface -----------------
--    GT0_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
--    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--    GT0_GTHTXN_OUT                          : out  std_logic;
--    GT0_GTHTXP_OUT                          : out  std_logic;
--    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--    GT0_TXOUTCLK_OUT                        : out  std_logic;
--    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
--    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
--    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--    GT0_TXRESETDONE_OUT                     : out  std_logic;
--   
--    --_________________________________________________________________________
--    --_________________________________________________________________________
--    --GT1  (X1Y5)
--    --____________________________CHANNEL PORTS________________________________
--    --------------------------------- CPLL Ports -------------------------------
--    GT1_CPLLFBCLKLOST_OUT                   : out  std_logic;
--    GT1_CPLLLOCK_OUT                        : out  std_logic;
--    GT1_CPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT1_CPLLRESET_IN                        : in   std_logic;
--    -------------------------- Channel - Clocking Ports ------------------------
--    GT1_GTREFCLK0_IN                        : in   std_logic;
--    ---------------------------- Channel - DRP Ports  --------------------------
--    GT1_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
--    GT1_DRPCLK_IN                           : in   std_logic;
--    GT1_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
--    GT1_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
--    GT1_DRPEN_IN                            : in   std_logic;
--    GT1_DRPRDY_OUT                          : out  std_logic;
--    GT1_DRPWE_IN                            : in   std_logic;
--    --------------------- RX Initialization and Reset Ports --------------------
--    GT1_RXUSERRDY_IN                        : in   std_logic;
--    -------------------------- RX Margin Analysis Ports ------------------------
--    GT1_EYESCANDATAERROR_OUT                : out  std_logic;
--    ------------------------- Receive Ports - CDR Ports ------------------------
--    GT1_RXCDRLOCK_OUT                       : out  std_logic;
--    --------------- Receive Ports - Comma Detection and Alignment --------------
--    GT1_RXSLIDE_IN                          : in   std_logic;
--    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--    GT1_RXUSRCLK_IN                         : in   std_logic;
--    GT1_RXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Receive Ports - FPGA RX interface Ports -----------------
--    GT1_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
--    ------------------------ Receive Ports - RX AFE Ports ----------------------
--    GT1_GTHRXN_IN                           : in   std_logic;
--    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--    GT1_RXPHMONITOR_OUT                     : out  std_logic_vector(4 downto 0);
--    GT1_RXPHSLIPMONITOR_OUT                 : out  std_logic_vector(4 downto 0);
--    --------------- Receive Ports - RX Fabric Output Control Ports -------------
--    GT1_RXOUTCLK_OUT                        : out  std_logic;
--    ------------- Receive Ports - RX Initialization and Reset Ports ------------
--    GT1_GTRXRESET_IN                        : in   std_logic;
--    ------------------------ Receive Ports -RX AFE Ports -----------------------
--    GT1_GTHRXP_IN                           : in   std_logic;
--    -------------- Receive Ports -RX Initialization and Reset Ports ------------
--    GT1_RXRESETDONE_OUT                     : out  std_logic;
--    --------------------- TX Initialization and Reset Ports --------------------
--    GT1_GTTXRESET_IN                        : in   std_logic;
--    GT1_TXUSERRDY_IN                        : in   std_logic;
--    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--    GT1_TXUSRCLK_IN                         : in   std_logic;
--    GT1_TXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Transmit Ports - TX Data Path interface -----------------
--    GT1_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
--    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--    GT1_GTHTXN_OUT                          : out  std_logic;
--    GT1_GTHTXP_OUT                          : out  std_logic;
--    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--    GT1_TXOUTCLK_OUT                        : out  std_logic;
--    GT1_TXOUTCLKFABRIC_OUT                  : out  std_logic;
--    GT1_TXOUTCLKPCS_OUT                     : out  std_logic;
--    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--    GT1_TXRESETDONE_OUT                     : out  std_logic;
--   
--    --_________________________________________________________________________
--    --_________________________________________________________________________
--    --GT2  (X1Y6)
--    --____________________________CHANNEL PORTS________________________________
--    --------------------------------- CPLL Ports -------------------------------
--    GT2_CPLLFBCLKLOST_OUT                   : out  std_logic;
--    GT2_CPLLLOCK_OUT                        : out  std_logic;
--    GT2_CPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT2_CPLLRESET_IN                        : in   std_logic;
--    -------------------------- Channel - Clocking Ports ------------------------
--    GT2_GTREFCLK0_IN                        : in   std_logic;
--    ---------------------------- Channel - DRP Ports  --------------------------
--    GT2_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
--    GT2_DRPCLK_IN                           : in   std_logic;
--    GT2_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
--    GT2_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
--    GT2_DRPEN_IN                            : in   std_logic;
--    GT2_DRPRDY_OUT                          : out  std_logic;
--    GT2_DRPWE_IN                            : in   std_logic;
--    --------------------- RX Initialization and Reset Ports --------------------
--    GT2_RXUSERRDY_IN                        : in   std_logic;
--    -------------------------- RX Margin Analysis Ports ------------------------
--    GT2_EYESCANDATAERROR_OUT                : out  std_logic;
--    ------------------------- Receive Ports - CDR Ports ------------------------
--    GT2_RXCDRLOCK_OUT                       : out  std_logic;
--    --------------- Receive Ports - Comma Detection and Alignment --------------
--    GT2_RXSLIDE_IN                          : in   std_logic;
--    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--    GT2_RXUSRCLK_IN                         : in   std_logic;
--    GT2_RXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Receive Ports - FPGA RX interface Ports -----------------
--    GT2_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
--    ------------------------ Receive Ports - RX AFE Ports ----------------------
--    GT2_GTHRXN_IN                           : in   std_logic;
--    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--    GT2_RXPHMONITOR_OUT                     : out  std_logic_vector(4 downto 0);
--    GT2_RXPHSLIPMONITOR_OUT                 : out  std_logic_vector(4 downto 0);
--    --------------- Receive Ports - RX Fabric Output Control Ports -------------
--    GT2_RXOUTCLK_OUT                        : out  std_logic;
--    ------------- Receive Ports - RX Initialization and Reset Ports ------------
--    GT2_GTRXRESET_IN                        : in   std_logic;
--    ------------------------ Receive Ports -RX AFE Ports -----------------------
--    GT2_GTHRXP_IN                           : in   std_logic;
--    -------------- Receive Ports -RX Initialization and Reset Ports ------------
--    GT2_RXRESETDONE_OUT                     : out  std_logic;
--    --------------------- TX Initialization and Reset Ports --------------------
--    GT2_GTTXRESET_IN                        : in   std_logic;
--    GT2_TXUSERRDY_IN                        : in   std_logic;
--    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--    GT2_TXUSRCLK_IN                         : in   std_logic;
--    GT2_TXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Transmit Ports - TX Data Path interface -----------------
--    GT2_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
--    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--    GT2_GTHTXN_OUT                          : out  std_logic;
--    GT2_GTHTXP_OUT                          : out  std_logic;
--    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--    GT2_TXOUTCLK_OUT                        : out  std_logic;
--    GT2_TXOUTCLKFABRIC_OUT                  : out  std_logic;
--    GT2_TXOUTCLKPCS_OUT                     : out  std_logic;
--    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--    GT2_TXRESETDONE_OUT                     : out  std_logic;
--   
--    --_________________________________________________________________________
--    --_________________________________________________________________________
--    --GT3  (X1Y7)
--    --____________________________CHANNEL PORTS________________________________
--    --------------------------------- CPLL Ports -------------------------------
--    GT3_CPLLFBCLKLOST_OUT                   : out  std_logic;
--    GT3_CPLLLOCK_OUT                        : out  std_logic;
--    GT3_CPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT3_CPLLRESET_IN                        : in   std_logic;
--    -------------------------- Channel - Clocking Ports ------------------------
--    GT3_GTREFCLK0_IN                        : in   std_logic;
--    ---------------------------- Channel - DRP Ports  --------------------------
--    GT3_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
--    GT3_DRPCLK_IN                           : in   std_logic;
--    GT3_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
--    GT3_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
--    GT3_DRPEN_IN                            : in   std_logic;
--    GT3_DRPRDY_OUT                          : out  std_logic;
--    GT3_DRPWE_IN                            : in   std_logic;
--    --------------------- RX Initialization and Reset Ports --------------------
--    GT3_RXUSERRDY_IN                        : in   std_logic;
--    -------------------------- RX Margin Analysis Ports ------------------------
--    GT3_EYESCANDATAERROR_OUT                : out  std_logic;
--    ------------------------- Receive Ports - CDR Ports ------------------------
--    GT3_RXCDRLOCK_OUT                       : out  std_logic;
--    --------------- Receive Ports - Comma Detection and Alignment --------------
--    GT3_RXSLIDE_IN                          : in   std_logic;
--    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
--    GT3_RXUSRCLK_IN                         : in   std_logic;
--    GT3_RXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Receive Ports - FPGA RX interface Ports -----------------
--    GT3_RXDATA_OUT                          : out  std_logic_vector(19 downto 0);
--    ------------------------ Receive Ports - RX AFE Ports ----------------------
--    GT3_GTHRXN_IN                           : in   std_logic;
--    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
--    GT3_RXPHMONITOR_OUT                     : out  std_logic_vector(4 downto 0);
--    GT3_RXPHSLIPMONITOR_OUT                 : out  std_logic_vector(4 downto 0);
--    --------------- Receive Ports - RX Fabric Output Control Ports -------------
--    GT3_RXOUTCLK_OUT                        : out  std_logic;
--    ------------- Receive Ports - RX Initialization and Reset Ports ------------
--    GT3_GTRXRESET_IN                        : in   std_logic;
--    ------------------------ Receive Ports -RX AFE Ports -----------------------
--    GT3_GTHRXP_IN                           : in   std_logic;
--    -------------- Receive Ports -RX Initialization and Reset Ports ------------
--    GT3_RXRESETDONE_OUT                     : out  std_logic;
--    --------------------- TX Initialization and Reset Ports --------------------
--    GT3_GTTXRESET_IN                        : in   std_logic;
--    GT3_TXUSERRDY_IN                        : in   std_logic;
--    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
--    GT3_TXUSRCLK_IN                         : in   std_logic;
--    GT3_TXUSRCLK2_IN                        : in   std_logic;
--    ------------------ Transmit Ports - TX Data Path interface -----------------
--    GT3_TXDATA_IN                           : in   std_logic_vector(19 downto 0);
--    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
--    GT3_GTHTXN_OUT                          : out  std_logic;
--    GT3_GTHTXP_OUT                          : out  std_logic;
--    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
--    GT3_TXOUTCLK_OUT                        : out  std_logic;
--    GT3_TXOUTCLKFABRIC_OUT                  : out  std_logic;
--    GT3_TXOUTCLKPCS_OUT                     : out  std_logic;
--    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
--    GT3_TXRESETDONE_OUT                     : out  std_logic;
--   
--
--    --____________________________COMMON PORTS________________________________
--    ---------------------- Common Block  - Ref Clock Ports ---------------------
--    GT0_GTREFCLK0_COMMON_IN                 : in   std_logic;
--    ------------------------- Common Block - QPLL Ports ------------------------
--    GT0_QPLLLOCK_OUT                        : out  std_logic;
--    GT0_QPLLLOCKDETCLK_IN                   : in   std_logic;
--    GT0_QPLLRESET_IN                        : in   std_logic
--
--
--);
--end component;
--

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

    signal   gt0_txfsmresetdone_i            : std_logic;
    signal   gt0_rxfsmresetdone_i            : std_logic;
    signal   gt0_txfsmresetdone_r            : std_logic;
    signal   gt0_txfsmresetdone_r2           : std_logic;
    signal   gt0_rxresetdone_r               : std_logic;
    signal   gt0_rxresetdone_r2              : std_logic;
    signal   gt0_rxresetdone_r3              : std_logic;


    signal   gt1_txfsmresetdone_i            : std_logic;
    signal   gt1_rxfsmresetdone_i            : std_logic;
    signal   gt1_txfsmresetdone_r            : std_logic;
    signal   gt1_txfsmresetdone_r2           : std_logic;
    signal   gt1_rxresetdone_r               : std_logic;
    signal   gt1_rxresetdone_r2              : std_logic;
    signal   gt1_rxresetdone_r3              : std_logic;


    signal   gt2_txfsmresetdone_i            : std_logic;
    signal   gt2_rxfsmresetdone_i            : std_logic;
    signal   gt2_txfsmresetdone_r            : std_logic;
    signal   gt2_txfsmresetdone_r2           : std_logic;
    signal   gt2_rxresetdone_r               : std_logic;
    signal   gt2_rxresetdone_r2              : std_logic;
    signal   gt2_rxresetdone_r3              : std_logic;


    signal   gt3_txfsmresetdone_i            : std_logic;
    signal   gt3_rxfsmresetdone_i            : std_logic;
    signal   gt3_txfsmresetdone_r            : std_logic;
    signal   gt3_txfsmresetdone_r2           : std_logic;
    signal   gt3_rxresetdone_r               : std_logic;
    signal   gt3_rxresetdone_r2              : std_logic;
    signal   gt3_rxresetdone_r3              : std_logic;



--**************************** Wire Declarations ******************************
    -------------------------- GT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GT0   (X1Y4)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt0_cpllfbclklost_out             : std_logic;
    signal  gt0_cplllock_out                  : std_logic;
    signal  gt0_cpllrefclklost_out            : std_logic;
    signal  gt0_cpllreset_in                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt0_drpaddr_in                   : std_logic_vector(8 downto 0);
    signal  gt0_drpdi_in                     : std_logic_vector(15 downto 0);
    signal  gt0_drpdo_out                     : std_logic_vector(15 downto 0);
    signal  gt0_drpen_in                     : std_logic;
    signal  gt0_drprdy_out                    : std_logic;
    signal  gt0_drpwe_in                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt0_rxuserrdy_in                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt0_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt0_rxcdrlock_i                 : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt0_rxslide_ni                   : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt0_rxdata_out                    : std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt0_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt0_rxdlyen_i                   : std_logic;
    signal  gt0_rxdlysreset_i               : std_logic;
    signal  gt0_rxdlysresetdone_i           : std_logic;
    signal  gt0_rxphalign_i                 : std_logic;
    signal  gt0_rxphaligndone_i             : std_logic;
    signal  gt0_rxphalignen_i               : std_logic;
    signal  gt0_rxphdlyreset_i              : std_logic;
    signal  gt0_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt0_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt0_rxsyncallin_i               : std_logic;
    signal  gt0_rxsyncdone_i                : std_logic;
    signal  gt0_rxsyncin_i                  : std_logic;
    signal  gt0_rxsyncmode_i                : std_logic;
    signal  gt0_rxsyncout_i                 : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt0_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt0_gtrxreset_iN                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt0_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt0_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt0_gttxreset_in                 : std_logic;
    signal  gt0_txuserrdy_in                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt0_txdlyen_i                   : std_logic;
    signal  gt0_txdlysreset_i               : std_logic;
    signal  gt0_txdlysresetdone_i           : std_logic;
    signal  gt0_txphalign_i                 : std_logic;
    signal  gt0_txphaligndone_i             : std_logic;
    signal  gt0_txphalignen_i               : std_logic;
    signal  gt0_txphdlyreset_i              : std_logic;
    signal  gt0_txphinit_i                  : std_logic;
    signal  gt0_txphinitdone_i              : std_logic;
    signal  gt0_txsyncallin_i               : std_logic;
    signal  gt0_txsyncdone_i                : std_logic;
    signal  gt0_txsyncin_i                  : std_logic;
    signal  gt0_txsyncmode_i                : std_logic;
    signal  gt0_txsyncout_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt0_txdata_in                    : std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt0_gthtxn_i                    : std_logic;
    signal  gt0_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt0_txoutclk_i                  : std_logic;
    signal  gt0_txoutclkfabric_i            : std_logic;
    signal  gt0_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt0_txresetdone_i               : std_logic;


    --________________________________________________________________________
    --________________________________________________________________________
    --GT1   (X1Y5)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt1_cpllfbclklost_out             : std_logic;
    signal  gt1_cplllock_out                  : std_logic;
    signal  gt1_cpllrefclklost_out            : std_logic;
    signal  gt1_cpllreset_in                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt1_drpaddr_in                   : std_logic_vector(8 downto 0);
    signal  gt1_drpdi_in                     : std_logic_vector(15 downto 0);
    signal  gt1_drpdo_out                     : std_logic_vector(15 downto 0);
    signal  gt1_drpen_in                     : std_logic;
    signal  gt1_drprdy_out                    : std_logic;
    signal  gt1_drpwe_in                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt1_rxuserrdy_in                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt1_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt1_rxcdrlock_i                 : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt1_rxslide_in                   : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt1_rxdata_OUT                    : std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt1_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt1_rxdlyen_i                   : std_logic;
    signal  gt1_rxdlysreset_i               : std_logic;
    signal  gt1_rxdlysresetdone_i           : std_logic;
    signal  gt1_rxphalign_i                 : std_logic;
    signal  gt1_rxphaligndone_i             : std_logic;
    signal  gt1_rxphalignen_i               : std_logic;
    signal  gt1_rxphdlyreset_i              : std_logic;
    signal  gt1_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt1_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt1_rxsyncallin_i               : std_logic;
    signal  gt1_rxsyncdone_i                : std_logic;
    signal  gt1_rxsyncin_i                  : std_logic;
    signal  gt1_rxsyncmode_i                : std_logic;
    signal  gt1_rxsyncout_i                 : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt1_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt1_gtrxreset_in                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt1_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt1_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt1_gttxreset_in                 : std_logic;
    signal  gt1_txuserrdy_in                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt1_txdlyen_i                   : std_logic;
    signal  gt1_txdlysreset_i               : std_logic;
    signal  gt1_txdlysresetdone_i           : std_logic;
    signal  gt1_txphalign_i                 : std_logic;
    signal  gt1_txphaligndone_i             : std_logic;
    signal  gt1_txphalignen_i               : std_logic;
    signal  gt1_txphdlyreset_i              : std_logic;
    signal  gt1_txphinit_i                  : std_logic;
    signal  gt1_txphinitdone_i              : std_logic;
    signal  gt1_txsyncallin_i               : std_logic;
    signal  gt1_txsyncdone_i                : std_logic;
    signal  gt1_txsyncin_i                  : std_logic;
    signal  gt1_txsyncmode_i                : std_logic;
    signal  gt1_txsyncout_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt1_txdata_in                    : std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt1_gthtxn_i                    : std_logic;
    signal  gt1_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt1_txoutclk_i                  : std_logic;
    signal  gt1_txoutclkfabric_i            : std_logic;
    signal  gt1_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt1_txresetdone_out               : std_logic;


    --________________________________________________________________________
    --________________________________________________________________________
    --GT2   (X1Y6)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt2_cpllfbclklost_out             : std_logic;
    signal  gt2_cplllock_out                  : std_logic;
    signal  gt2_cpllrefclklost_out            : std_logic;
    signal  gt2_cpllreset_in                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt2_drpaddr_in                   : std_logic_vector(8 downto 0);
    signal  gt2_drpdi_in                     : std_logic_vector(15 downto 0);
    signal  gt2_drpdo_out                     : std_logic_vector(15 downto 0);
    signal  gt2_drpen_in                     : std_logic;
    signal  gt2_drprdy_out                    : std_logic;
    signal  gt2_drpwe_in                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt2_rxuserrdy_in                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt2_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt2_rxcdrlock_i                 : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt2_rxslide_in                   : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt2_rxdata_OUT                    : std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt2_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt2_rxdlyen_i                   : std_logic;
    signal  gt2_rxdlysreset_i               : std_logic;
    signal  gt2_rxdlysresetdone_i           : std_logic;
    signal  gt2_rxphalign_i                 : std_logic;
    signal  gt2_rxphaligndone_i             : std_logic;
    signal  gt2_rxphalignen_i               : std_logic;
    signal  gt2_rxphdlyreset_i              : std_logic;
    signal  gt2_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt2_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt2_rxsyncallin_i               : std_logic;
    signal  gt2_rxsyncdone_i                : std_logic;
    signal  gt2_rxsyncin_i                  : std_logic;
    signal  gt2_rxsyncmode_i                : std_logic;
    signal  gt2_rxsyncout_i                 : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt2_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt2_gtrxreset_in                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt2_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt2_rxresetdone_out               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt2_gttxreset_in                 : std_logic;
    signal  gt2_txuserrdy_in                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt2_txdlyen_i                   : std_logic;
    signal  gt2_txdlysreset_i               : std_logic;
    signal  gt2_txdlysresetdone_i           : std_logic;
    signal  gt2_txphalign_i                 : std_logic;
    signal  gt2_txphaligndone_i             : std_logic;
    signal  gt2_txphalignen_i               : std_logic;
    signal  gt2_txphdlyreset_i              : std_logic;
    signal  gt2_txphinit_i                  : std_logic;
    signal  gt2_txphinitdone_i              : std_logic;
    signal  gt2_txsyncallin_i               : std_logic;
    signal  gt2_txsyncdone_i                : std_logic;
    signal  gt2_txsyncin_i                  : std_logic;
    signal  gt2_txsyncmode_i                : std_logic;
    signal  gt2_txsyncout_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt2_txdata_in                    : std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt2_gthtxn_i                    : std_logic;
    signal  gt2_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt2_txoutclk_i                  : std_logic;
    signal  gt2_txoutclkfabric_i            : std_logic;
    signal  gt2_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt2_txresetdone_i               : std_logic;


    --________________________________________________________________________
    --________________________________________________________________________
    --GT3   (X1Y7)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt3_cpllfbclklost_out             : std_logic;
    signal  gt3_cplllock_out                  : std_logic;
    signal  gt3_cpllrefclklost_out            : std_logic;
    signal  gt3_cpllreset_in                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt3_drpaddr_iN                   : std_logic_vector(8 downto 0);
    signal  gt3_drpdi_iN                     : std_logic_vector(15 downto 0);
    signal  gt3_drpdo_out                     : std_logic_vector(15 downto 0);
    signal  gt3_drpen_in                     : std_logic;
    signal  gt3_drprdy_out                    : std_logic;
    signal  gt3_drpwe_in                     : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt3_rxuserrdy_ni                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt3_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt3_rxcdrlock_i                 : std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  gt3_rxslide_in                   : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt3_rxdata_OUT                    : std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt3_gthrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt3_rxdlyen_i                   : std_logic;
    signal  gt3_rxdlysreset_i               : std_logic;
    signal  gt3_rxdlysresetdone_i           : std_logic;
    signal  gt3_rxphalign_i                 : std_logic;
    signal  gt3_rxphaligndone_i             : std_logic;
    signal  gt3_rxphalignen_i               : std_logic;
    signal  gt3_rxphdlyreset_i              : std_logic;
    signal  gt3_rxphmonitor_i               : std_logic_vector(4 downto 0);
    signal  gt3_rxphslipmonitor_i           : std_logic_vector(4 downto 0);
    signal  gt3_rxsyncallin_i               : std_logic;
    signal  gt3_rxsyncdone_i                : std_logic;
    signal  gt3_rxsyncin_i                  : std_logic;
    signal  gt3_rxsyncmode_i                : std_logic;
    signal  gt3_rxsyncout_i                 : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt3_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt3_gtrxreset_in                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt3_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt3_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt3_gttxreset_in                 : std_logic;
    signal  gt3_txuserrdy_in                 : std_logic;
    ------------------ Transmit Ports - TX Buffer Bypass Ports -----------------
    signal  gt3_txdlyen_i                   : std_logic;
    signal  gt3_txdlysreset_i               : std_logic;
    signal  gt3_txdlysresetdone_i           : std_logic;
    signal  gt3_txphalign_i                 : std_logic;
    signal  gt3_txphaligndone_i             : std_logic;
    signal  gt3_txphalignen_i               : std_logic;
    signal  gt3_txphdlyreset_i              : std_logic;
    signal  gt3_txphinit_i                  : std_logic;
    signal  gt3_txphinitdone_i              : std_logic;
    signal  gt3_txsyncallin_i               : std_logic;
    signal  gt3_txsyncdone_i                : std_logic;
    signal  gt3_txsyncin_i                  : std_logic;
    signal  gt3_txsyncmode_i                : std_logic;
    signal  gt3_txsyncout_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt3_txdata_iN                    : std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt3_gthtxn_i                    : std_logic;
    signal  gt3_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt3_txoutclk_i                  : std_logic;
    signal  gt3_txoutclkfabric_i            : std_logic;
    signal  gt3_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt3_txresetdone_i               : std_logic;



    --____________________________COMMON PORTS________________________________
    ------------------------- Common Block - QPLL Ports ------------------------
    signal  gt0_qplllock_i                  : std_logic;
    signal  gt0_qpllrefclklost_i            : std_logic;
    signal  gt0_qpllreset_i                 : std_logic;



    ------------------------------- Global Signals -----------------------------
    signal  gt0_tx_system_reset_c           : std_logic;
    signal  gt0_rx_system_reset_c           : std_logic;
    signal  gt1_tx_system_reset_c           : std_logic;
    signal  gt1_rx_system_reset_c           : std_logic;
    signal  gt2_tx_system_reset_c           : std_logic;
    signal  gt2_rx_system_reset_c           : std_logic;
    signal  gt3_tx_system_reset_c           : std_logic;
    signal  gt3_rx_system_reset_c           : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drpclk_in_i                     : std_logic;
 
    signal  GTTXRESET_IN                    : std_logic;
    signal  GTRXRESET_IN                    : std_logic;
    signal  CPLLRESET_IN                    : std_logic;
    signal  QPLLRESET_IN                    : std_logic;

   ------------------------------- User Clocks ---------------------------------
    attribute keep: string;
  --  signal    gt0_txusrclk_in                  : std_logic; 
    signal    gt0_txusrclk2_in                 : std_logic; 
  --  signal    gt0_rxusrclk_i                  : std_logic; 
    signal    gt0_rxusrclk2_in                 : std_logic; 
    attribute keep of gt0_txusrclk_in : signal is "true";
    attribute keep of gt0_txusrclk2_in : signal is "true";
    --attribute keep of gt0_rxusrclk_i : signal is "true";
    attribute keep of gt0_rxusrclk2_in : signal is "true";
   signal    gt1_txusrclk_in                  : std_logic; 
    signal    gt1_txusrclk2_in                 : std_logic; 
  --  signal    gt1_rxusrclk_i                  : std_logic; 
    signal    gt1_rxusrclk2_in                 : std_logic; 
    attribute keep of gt1_txusrclk_in : signal is "true";
    attribute keep of gt1_txusrclk2_in : signal is "true";
  --  attribute keep of gt1_rxusrclk_in : signal is "true";
    attribute keep of gt1_rxusrclk2_in : signal is "true";
    signal    gt2_txusrclk_in                  : std_logic; 
    signal    gt2_txusrclk2_in                 : std_logic; 
   -- signal    gt2_rxusrclk_in                  : std_logic; 
    signal    gt2_rxusrclk2_in                 : std_logic; 
    attribute keep of gt2_txusrclk_in : signal is "true";
    attribute keep of gt2_txusrclk2_in : signal is "true";
   -- attribute keep of gt2_rxusrclk_i : signal is "true";
    attribute keep of gt2_rxusrclk2_in : signal is "true";
    signal    gt3_txusrclk_in                  : std_logic; 
    signal    gt3_txusrclk2_in                 : std_logic; 
   -- signal    gt3_rxusrclk_in                  : std_logic; 
    signal    gt3_rxusrclk2_in                 : std_logic; 
    attribute keep of gt3_txusrclk_in : signal is "true";
    attribute keep of gt3_txusrclk2_in : signal is "true";
   -- attribute keep of gt3_rxusrclk_i : signal is "true";
    attribute keep of gt3_rxusrclk2_in : signal is "true";
 

signal gt2_txoutclk_out,gt1_txoutclk_out, gt3_txoutclk_out:std_logic;

    ----------------------------- Reference Clocks ----------------------------
    signal gt3_rxuserrdy_in:std_logic;
    signal    q2_clk0_refclk_i                : std_logic;

signal GT0_TX_FSM_RESET_DONE_OUT,GT1_TX_FSM_RESET_DONE_OUT,GT2_TX_FSM_RESET_DONE_OUT,GT3_TX_FSM_RESET_DONE_OUT:std_logic;
signal GT0_RX_FSM_RESET_DONE_OUT,GT1_RX_FSM_RESET_DONE_OUT,GT2_RX_FSM_RESET_DONE_OUT,GT3_RX_FSM_RESET_DONE_OUT:std_logic;
   signal gt0_gtrefclk0_in,gt1_gtrefclk0_in,gt2_gtrefclk0_in,gt3_gtrefclk0_in,gt3_rxresetdone_out,gt1_rxresetdone_out: std_logic;
signal gt3_txresetdone_out,gt2_txresetdone_out,gt0_txresetdone_out,gt0_rxslide_in,gt0_rxresetdone_out:std_logic;
--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_ground_vec_i                         <= x"0000000000000000";
    tied_to_vcc_i                                <= '1';
    tied_to_vcc_vec_i                            <= x"ff";

----------------------------
------- edited by C.K.   
    --CONNECTIONs added
	 drpclk_in_i 		<= 	DRP_CLK_IN;
	 --q2_clk0_refclk_i <= 	q2_clk0_refclk_in; 
	 gt1_gtrefclk0_in<= 	q2_clk0_refclk_in; 
	  gt2_gtrefclk0_in<= 	q2_clk0_refclk_in; 
	   gt3_gtrefclk0_in<= 	q2_clk0_refclk_in; 
	    gt0_gtrefclk0_in<= 	q2_clk0_refclk_in; 
	 gt3_rxslide_in <= gt_rxslide_in(3);
	 gt2_rxslide_in <= gt_rxslide_in(2);
	 gt1_rxslide_in <= gt_rxslide_in(1);
	 gt0_rxslide_in <= gt_rxslide_in(0);
	 
	 gt0_txuserrdy_in <= gt_txuserrdy_in(0);
	 gt1_txuserrdy_in <= gt_txuserrdy_in(1);
	 gt2_txuserrdy_in <= gt_txuserrdy_in(2);
	 gt3_txuserrdy_in <= gt_txuserrdy_in(3);
	  gt0_rxuserrdy_in <= gt_rxuserrdy_in(0);
         gt1_rxuserrdy_in <= gt_rxuserrdy_in(1);
         gt2_rxuserrdy_in <= gt_rxuserrdy_in(2);
         gt3_rxuserrdy_in <= gt_rxuserrdy_in(3);
	 
	 gt0_qpllreset_i <= QPLL_RESET_IN;
	 
	 gt0_cpllreset_in <= CPLL_RESET_IN(0);
	 gt1_cpllreset_in <= CPLL_RESET_IN(1);
	 gt2_cpllreset_in <= CPLL_RESET_IN(2);
	 gt3_cpllreset_in <= CPLL_RESET_IN(3);
	 
	 gt0_gtrxreset_in                              <= GTRX_RESET_IN(0) or not gt0_cplllock_OUT;
    gt0_gttxreset_in                              <= GTTX_RESET_IN(0) or not gt0_cplllock_OUT;
	 gt1_gtrxreset_in                              <= GTRX_RESET_IN(1) or not gt1_cplllock_OUT;
    gt1_gttxreset_in                              <= GTTX_RESET_IN(1) or not gt1_cplllock_OUT;
	 gt2_gtrxreset_in                              <= GTRX_RESET_IN(2) or not gt2_cplllock_OUT;
    gt2_gttxreset_in                              <= GTTX_RESET_IN(2) or not gt2_cplllock_OUT;
	 gt3_gtrxreset_in                              <= GTRX_RESET_IN(3) or not gt3_cplllock_OUT;
    gt3_gttxreset_in                              <= GTTX_RESET_IN(3) or not gt3_cplllock_OUT;
    
  
	 gt_txfsmresetdone_out 	<= 	GT3_TX_FSM_RESET_DONE_OUT & GT2_TX_FSM_RESET_DONE_OUT & GT1_TX_FSM_RESET_DONE_OUT & GT0_TX_FSM_RESET_DONE_OUT;
	 gt_rxfsmresetdone_out 	<= GT3_RX_FSM_RESET_DONE_OUT & GT2_RX_FSM_RESET_DONE_OUT & GT1_RX_FSM_RESET_DONE_OUT & GT0_RX_FSM_RESET_DONE_OUT;
	 
	 gt_txresetdone_out    	<= 	gt3_txresetdone_out & gt2_txresetdone_out & gt1_txresetdone_out & gt0_txresetdone_out;
	 gt_rxresetdone_out    	<= 	gt3_rxresetdone_out & gt2_rxresetdone_out & gt1_rxresetdone_out & gt0_rxresetdone_out;
	 
	 gt_cpllfbclklost_out 	<= 	gt3_cpllfbclklost_out & gt2_cpllfbclklost_out & gt1_cpllfbclklost_out & gt0_cpllfbclklost_out;
	 gt_cplllock_OUT 			<= 	gt3_cplllock_out & gt2_cplllock_out & gt1_cplllock_out & gt0_cplllock_out;
	 gt_rxcdrlock_OUT 		<= 	"1111";--gt3_rxcdrlock_i & gt2_rxcdrlock_i & gt1_rxcdrlock_i & gt0_rxcdrlock_i;
	 
	 gt_qplllock_out <= gt0_qplllock_i;
	 
	 
	 gt0_txdata_in <= TX_DATA_gt0_20b;
	 gt1_txdata_in <= TX_DATA_gt1_20b;
	 gt2_txdata_in <= TX_DATA_gt2_20b;
	 gt3_txdata_in <= TX_DATA_gt3_20b;
	 RX_DATA_gt0_20b <= gt0_rxdata_out;
	 RX_DATA_gt1_20b <= gt1_rxdata_out;
	 RX_DATA_gt2_20b <= gt2_rxdata_out;
	 RX_DATA_gt3_20b <= gt3_rxdata_out;
	 
	 
	 gt0_rxusrclk2_in 	<= gt0_rxusrclk_in;
	-- gt0_rxusrclk_in 	<= gt0_rxusrclk_in;
	-- gt0_rxoutclk_out <= gt0_rxoutclk_out;
	 
	 gt1_rxusrclk2_in 	<= gt1_rxusrclk_in;
	-- gt1_rxusrclk_in 	<= gt1_rxusrclk_in;
	-- gt1_rxoutclk_out <= gt1_rxoutclk_out;
	 
	 gt2_rxusrclk2_in 	<= gt2_rxusrclk_in;
	 --gt2_rxusrclk_in 	<= gt2_rxusrclk_in;
--	 gt2_rxoutclk_out <= gt2_rxoutclk_out;
	 
	 gt3_rxusrclk2_in 	<= gt3_rxusrclk_in;
	 --gt3_rxusrclk_in 	<= gt3_rxusrclk_in;
--	 gt3_rxoutclk_out <= gt3_rxoutclk_out;
	 
	 gt0_txusrclk2_in 	<= gt0_txusrclk_in;
	-- gt0_txusrclk_in 	<= gt0_txusrclk_in;
	-- gt0_txoutclk_out <= gt0_txoutclk_out;
	 
	 gt1_txusrclk2_in 	<= gt0_txusrclk_in;
	 gt1_txusrclk_in 	<= gt0_txusrclk_in;
	 gt2_txusrclk2_in 	<= gt0_txusrclk_in;
	 gt2_txusrclk_in 	<= gt0_txusrclk_in;
	 gt3_txusrclk2_in 	<= gt0_txusrclk_in;
	 gt3_txusrclk_in 	<= gt0_txusrclk_in;
	 
    
  
  
      gth_quad_4p8g_cpll_init_i : entity work.gth_quad_4p8g_cpll_manual_init
      generic map
  (
          EXAMPLE_SIM_GTRESET_SPEEDUP   => "TRUE",
          EXAMPLE_SIMULATION            => 0,
   
          STABLE_CLOCK_PERIOD           => STABLE_CLOCK_PERIOD,
          EXAMPLE_USE_CHIPSCOPE         => 1
  )
  port map
  (
          SYSCLK_IN                       =>     drpclk_in_i,-- SYSCLK_IN,
          SOFT_RESET_IN                   =>      SOFT_RESET_IN,
           SOFT_TXRST_GT       =>  SOFT_TXRST_GT,
             SOFT_RXRST_GT       =>  SOFT_RXRST_GT,
             SOFT_TXRST_ALL      => SOFT_TXRST_ALL,
             SOFT_RXRST_ALL      => SOFT_RXRST_ALL,
          DONT_RESET_ON_DATA_ERROR_IN     =>     '1',-- DONT_RESET_ON_DATA_ERROR_IN,
      GT0_TX_FSM_RESET_DONE_OUT => GT0_TX_FSM_RESET_DONE_OUT,
      GT0_RX_FSM_RESET_DONE_OUT => GT0_RX_FSM_RESET_DONE_OUT,
      GT0_DATA_VALID_IN => '1',--GT0_DATA_VALID_IN,
      GT1_TX_FSM_RESET_DONE_OUT => GT1_TX_FSM_RESET_DONE_OUT,
      GT1_RX_FSM_RESET_DONE_OUT => GT1_RX_FSM_RESET_DONE_OUT,
      GT1_DATA_VALID_IN =>'1',-- GT1_DATA_VALID_IN,
      GT2_TX_FSM_RESET_DONE_OUT => GT2_TX_FSM_RESET_DONE_OUT,
      GT2_RX_FSM_RESET_DONE_OUT => GT2_RX_FSM_RESET_DONE_OUT,
      GT2_DATA_VALID_IN => '1',--GT2_DATA_VALID_IN,
      GT3_TX_FSM_RESET_DONE_OUT => GT3_TX_FSM_RESET_DONE_OUT,
      GT3_RX_FSM_RESET_DONE_OUT => GT3_RX_FSM_RESET_DONE_OUT,
      GT3_DATA_VALID_IN => '1',--GT3_DATA_VALID_IN,
  
      --_________________________________________________________________________
      --GT0  (X1Y4)
      --____________________________CHANNEL PORTS________________________________
      --------------------------------- CPLL Ports -------------------------------
          gt0_cpllfbclklost_out           =>      gt0_cpllfbclklost_out,
          gt0_cplllock_out                =>      gt0_cplllock_out,
          gt0_cplllockdetclk_in           =>       drpclk_in_i,--gt0_cplllockdetclk_in,
          gt0_cpllreset_in                =>      gt0_cpllreset_in,
      -------------------------- Channel - Clocking Ports ------------------------
          gt0_gtrefclk0_in                =>     gt0_gtrefclk0_in,
      ---------------------------- Channel - DRP Ports  --------------------------
          gt0_drpaddr_in                  =>      gt0_drpaddr_in,
          gt0_drpclk_in                   =>       drpclk_in_i,--gt0_drpclk_in,
          gt0_drpdi_in                    =>      gt0_drpdi_in,
          gt0_drpdo_out                   =>      gt0_drpdo_out,
          gt0_drpen_in                    =>      gt0_drpen_in,
          gt0_drprdy_out                  =>      open,--gt0_drprdy_out,
          gt0_drpwe_in                    =>      gt0_drpwe_in,
      --------------------- RX Initialization and Reset Ports --------------------
          gt0_eyescanreset_in             =>      '0',--gt0_eyescanreset_in,
          gt0_rxuserrdy_in                =>      gt0_rxuserrdy_in,
      -------------------------- RX Margin Analysis Ports ------------------------
          gt0_eyescandataerror_out        =>      open,--gt0_eyescandataerror_out,
          gt0_eyescantrigger_in           =>      '0',--gt0_eyescantrigger_in,
      --------------- Receive Ports - Comma Detection and Alignment --------------
          gt0_rxslide_in                  =>      gt0_rxslide_in,
      ------------------- Receive Ports - Digital Monitor Ports ------------------
          gt0_dmonitorout_out             =>    open,--  gt0_dmonitorout_out,
      ------------------ Receive Ports - FPGA RX Interface Ports -----------------
          gt0_rxusrclk_in                 =>      gt0_rxusrclk_in,
          gt0_rxusrclk2_in                =>      gt0_rxusrclk2_in,
      ------------------ Receive Ports - FPGA RX interface Ports -----------------
          gt0_rxdata_out                  =>      gt0_rxdata_out,
      ------------------------ Receive Ports - RX AFE Ports ----------------------
          gt0_gthrxn_in                   =>      RXN_IN(0),--gt0_gthrxn_in,
      ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
          gt0_rxphmonitor_out             =>   open,--    gt0_rxphmonitor_out,
          gt0_rxphslipmonitor_out         =>    open,--   gt0_rxphslipmonitor_out,
      --------------------- Receive Ports - RX Equalizer Ports -------------------
          gt0_rxmonitorout_out            =>   open,--    gt0_rxmonitorout_out,
          gt0_rxmonitorsel_in             =>   "00",--   gt0_rxmonitorsel_in,
      --------------- Receive Ports - RX Fabric Output Control Ports -------------
          gt0_rxoutclk_out                =>      gt0_rxoutclk_out,
      ------------- Receive Ports - RX Initialization and Reset Ports ------------
          gt0_gtrxreset_in                =>      gt0_gtrxreset_in,
      ------------------------ Receive Ports -RX AFE Ports -----------------------
          gt0_gthrxp_in                   =>        RXP_IN(0),--gt0_gthrxp_in,
      -------------- Receive Ports -RX Initialization and Reset Ports ------------
          gt0_rxresetdone_out             =>      gt0_rxresetdone_out,
      --------------------- TX Initialization and Reset Ports --------------------
          gt0_gttxreset_in                =>      gt0_gttxreset_in,
          gt0_txuserrdy_in                =>      gt0_txuserrdy_in,
      ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
          gt0_txusrclk_in                 =>      gt0_txusrclk_in,
          gt0_txusrclk2_in                =>      gt0_txusrclk2_in,
      ------------------ Transmit Ports - TX Data Path interface -----------------
          gt0_txdata_in                   =>      gt0_txdata_in,
      ---------------- Transmit Ports - TX Driver and OOB signaling --------------
          gt0_gthtxn_out                  =>        TXN_OUT(0),--gt0_gthtxn_out,
          gt0_gthtxp_out                  =>       TXP_OUT(0),-- gt0_gthtxp_out,
      ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
          gt0_txoutclk_out                =>      gt0_txoutclk_out,
          gt0_txoutclkfabric_out          =>      open,--gt0_txoutclkfabric_out,
          gt0_txoutclkpcs_out             =>      open,--gt0_txoutclkpcs_out,
      ------------- Transmit Ports - TX Initialization and Reset Ports -----------
          gt0_txresetdone_out             =>      gt0_txresetdone_out,
  
      --GT1  (X1Y5)
      --____________________________CHANNEL PORTS________________________________
      --------------------------------- CPLL Ports -------------------------------
          gt1_cpllfbclklost_out           =>      gt1_cpllfbclklost_out,
          gt1_cplllock_out                =>      gt1_cplllock_out,
          gt1_cplllockdetclk_in           =>      drpclk_in_i,-- gt1_cplllockdetclk_in,
          gt1_cpllreset_in                =>      gt1_cpllreset_in,
      -------------------------- Channel - Clocking Ports ------------------------
          gt1_gtrefclk0_in                =>      gt1_gtrefclk0_in,
      ---------------------------- Channel - DRP Ports  --------------------------
          gt1_drpaddr_in                  =>      gt1_drpaddr_in,
          gt1_drpclk_in                   =>      drpclk_in_i,-- gt1_drpclk_in,
          gt1_drpdi_in                    =>      gt1_drpdi_in,
          gt1_drpdo_out                   =>      gt1_drpdo_out,
          gt1_drpen_in                    =>      gt1_drpen_in,
          gt1_drprdy_out                  =>      gt1_drprdy_out,
          gt1_drpwe_in                    =>      gt1_drpwe_in,
      --------------------- RX Initialization and Reset Ports --------------------
          gt1_eyescanreset_in             =>    '0',--  gt1_eyescanreset_in,
          gt1_rxuserrdy_in                =>      gt1_rxuserrdy_in,
      -------------------------- RX Margin Analysis Ports ------------------------
          gt1_eyescandataerror_out        =>      open,--gt1_eyescandataerror_out,
          gt1_eyescantrigger_in           =>    '0',--  gt1_eyescantrigger_in,
      --------------- Receive Ports - Comma Detection and Alignment --------------
          gt1_rxslide_in                  =>      gt1_rxslide_in,
      ------------------- Receive Ports - Digital Monitor Ports ------------------
          gt1_dmonitorout_out             =>     open,-- gt1_dmonitorout_out,
      ------------------ Receive Ports - FPGA RX Interface Ports -----------------
          gt1_rxusrclk_in                 =>      gt1_rxusrclk_in,
          gt1_rxusrclk2_in                =>      gt1_rxusrclk2_in,
      ------------------ Receive Ports - FPGA RX interface Ports -----------------
          gt1_rxdata_out                  =>      gt1_rxdata_out,
      ------------------------ Receive Ports - RX AFE Ports ----------------------
          gt1_gthrxn_in                   =>      RXN_IN(1),--gt1_gthrxn_in,
      ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
          gt1_rxphmonitor_out             =>   open,--    gt1_rxphmonitor_out,
          gt1_rxphslipmonitor_out         =>   open,--    gt1_rxphslipmonitor_out,
      --------------------- Receive Ports - RX Equalizer Ports -------------------
          gt1_rxmonitorout_out            =>   open,--    gt1_rxmonitorout_out,
          gt1_rxmonitorsel_in             =>    "00",----  gt1_rxmonitorsel_in,
      --------------- Receive Ports - RX Fabric Output Control Ports -------------
          gt1_rxoutclk_out                =>      gt1_rxoutclk_out,
      ------------- Receive Ports - RX Initialization and Reset Ports ------------
          gt1_gtrxreset_in                =>      gt1_gtrxreset_in,
      ------------------------ Receive Ports -RX AFE Ports -----------------------
          gt1_gthrxp_in                   =>      RXP_IN(1),--gt1_gthrxp_in,
      -------------- Receive Ports -RX Initialization and Reset Ports ------------
          gt1_rxresetdone_out             =>      gt1_rxresetdone_out,
      --------------------- TX Initialization and Reset Ports --------------------
          gt1_gttxreset_in                =>      gt1_gttxreset_in,
          gt1_txuserrdy_in                =>      gt1_txuserrdy_in,
      ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
          gt1_txusrclk_in                 =>      gt1_txusrclk_in,
          gt1_txusrclk2_in                =>      gt1_txusrclk2_in,
      ------------------ Transmit Ports - TX Data Path interface -----------------
          gt1_txdata_in                   =>      gt1_txdata_in,
      ---------------- Transmit Ports - TX Driver and OOB signaling --------------
          gt1_gthtxn_out                  =>     TXN_OUT(1),-- gt1_gthtxn_out,
          gt1_gthtxp_out                  =>     TXP_OUT(1),-- gt1_gthtxp_out,
      ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
          gt1_txoutclk_out                =>      gt1_txoutclk_out,
          gt1_txoutclkfabric_out          =>     open,-- gt1_txoutclkfabric_out,
          gt1_txoutclkpcs_out             =>      open,--  gt1_txoutclkpcs_out,
      ------------- Transmit Ports - TX Initialization and Reset Ports -----------
          gt1_txresetdone_out             =>      gt1_txresetdone_out,
  
      --GT2  (X1Y6)
      --____________________________CHANNEL PORTS________________________________
      --------------------------------- CPLL Ports -------------------------------
          gt2_cpllfbclklost_out           =>      gt2_cpllfbclklost_out,
          gt2_cplllock_out                =>      gt2_cplllock_out,
          gt2_cplllockdetclk_in           =>      drpclk_in_i,-- gt2_cplllockdetclk_in,
          gt2_cpllreset_in                =>      gt2_cpllreset_in,
      -------------------------- Channel - Clocking Ports ------------------------
          gt2_gtrefclk0_in                =>      gt2_gtrefclk0_in,
      ---------------------------- Channel - DRP Ports  --------------------------
          gt2_drpaddr_in                  =>      gt2_drpaddr_in,
          gt2_drpclk_in                   =>      drpclk_in_i,-- gt2_drpclk_in,
          gt2_drpdi_in                    =>      gt2_drpdi_in,
          gt2_drpdo_out                   =>      gt2_drpdo_out,
          gt2_drpen_in                    =>      gt2_drpen_in,
          gt2_drprdy_out                  =>      gt2_drprdy_out,
          gt2_drpwe_in                    =>      gt2_drpwe_in,
      --------------------- RX Initialization and Reset Ports --------------------
          gt2_eyescanreset_in             =>    '0',--  gt2_eyescanreset_in,
          gt2_rxuserrdy_in                =>      gt2_rxuserrdy_in,
      -------------------------- RX Margin Analysis Ports ------------------------
          gt2_eyescandataerror_out        =>    open,--  gt2_eyescandataerror_out,
          gt2_eyescantrigger_in           =>    '0',--  gt2_eyescantrigger_in,
      --------------- Receive Ports - Comma Detection and Alignment --------------
          gt2_rxslide_in                  =>      gt2_rxslide_in,
      ------------------- Receive Ports - Digital Monitor Ports ------------------
          gt2_dmonitorout_out             =>    open,--  gt2_dmonitorout_out,
      ------------------ Receive Ports - FPGA RX Interface Ports -----------------
          gt2_rxusrclk_in                 =>      gt2_rxusrclk_in,
          gt2_rxusrclk2_in                =>      gt2_rxusrclk2_in,
      ------------------ Receive Ports - FPGA RX interface Ports -----------------
          gt2_rxdata_out                  =>      gt2_rxdata_out,
      ------------------------ Receive Ports - RX AFE Ports ----------------------
          gt2_gthrxn_in                   =>     RXN_IN(2),-- gt2_gthrxn_in,
      ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
          gt2_rxphmonitor_out             =>   open,--    gt2_rxphmonitor_out,
          gt2_rxphslipmonitor_out         =>   open,--    gt2_rxphslipmonitor_out,
      --------------------- Receive Ports - RX Equalizer Ports -------------------
          gt2_rxmonitorout_out            =>  open,--     gt2_rxmonitorout_out,
          gt2_rxmonitorsel_in             =>   "00",----    gt2_rxmonitorsel_in,
      --------------- Receive Ports - RX Fabric Output Control Ports -------------
          gt2_rxoutclk_out                =>      gt2_rxoutclk_out,
      ------------- Receive Ports - RX Initialization and Reset Ports ------------
          gt2_gtrxreset_in                =>      gt2_gtrxreset_in,
      ------------------------ Receive Ports -RX AFE Ports -----------------------
          gt2_gthrxp_in                   =>      RXP_IN(2),-- gt2_gthrxp_in,
      -------------- Receive Ports -RX Initialization and Reset Ports ------------
          gt2_rxresetdone_out             =>      gt2_rxresetdone_out,
      --------------------- TX Initialization and Reset Ports --------------------
          gt2_gttxreset_in                =>      gt2_gttxreset_in,
          gt2_txuserrdy_in                =>      gt2_txuserrdy_in,
      ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
          gt2_txusrclk_in                 =>      gt2_txusrclk_in,
          gt2_txusrclk2_in                =>      gt2_txusrclk2_in,
      ------------------ Transmit Ports - TX Data Path interface -----------------
          gt2_txdata_in                   =>      gt2_txdata_in,
      ---------------- Transmit Ports - TX Driver and OOB signaling --------------
          gt2_gthtxn_out                  =>     TXN_OUT(2),-- gt1_gthtxn_out,
                gt2_gthtxp_out                  =>     TXP_OUT(2),-- gt1_gthtxp_out,
      ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
          gt2_txoutclk_out                =>      gt2_txoutclk_out,
          gt2_txoutclkfabric_out          =>       open,-- gt2_txoutclkfabric_out,
          gt2_txoutclkpcs_out             =>      open,--  gt2_txoutclkpcs_out,
      ------------- Transmit Ports - TX Initialization and Reset Ports -----------
          gt2_txresetdone_out             =>      gt2_txresetdone_out,
  
      --GT3  (X1Y7)
      --____________________________CHANNEL PORTS________________________________
      --------------------------------- CPLL Ports -------------------------------
          gt3_cpllfbclklost_out           =>      gt3_cpllfbclklost_out,
          gt3_cplllock_out                =>      gt3_cplllock_out,
          gt3_cplllockdetclk_in           =>      drpclk_in_i,-- gt3_cplllockdetclk_in,
          gt3_cpllreset_in                =>      gt3_cpllreset_in,
      -------------------------- Channel - Clocking Ports ------------------------
          gt3_gtrefclk0_in                =>      gt3_gtrefclk0_in,
      ---------------------------- Channel - DRP Ports  --------------------------
          gt3_drpaddr_in                  =>      gt3_drpaddr_in,
          gt3_drpclk_in                   =>      drpclk_in_i,-- gt3_drpclk_in,
          gt3_drpdi_in                    =>      gt3_drpdi_in,
          gt3_drpdo_out                   =>      gt3_drpdo_out,
          gt3_drpen_in                    =>      gt3_drpen_in,
          gt3_drprdy_out                  =>      gt3_drprdy_out,
          gt3_drpwe_in                    =>      gt3_drpwe_in,
      --------------------- RX Initialization and Reset Ports --------------------
          gt3_eyescanreset_in             =>     '0',-- gt3_eyescanreset_in,
          gt3_rxuserrdy_in                =>      gt3_rxuserrdy_in,
      -------------------------- RX Margin Analysis Ports ------------------------
          gt3_eyescandataerror_out        =>   open,--   gt3_eyescandataerror_out,
          gt3_eyescantrigger_in           =>  '0',----   gt3_eyescantrigger_in,
      --------------- Receive Ports - Comma Detection and Alignment --------------
          gt3_rxslide_in                  =>      gt3_rxslide_in,
      ------------------- Receive Ports - Digital Monitor Ports ------------------
          gt3_dmonitorout_out             =>     open,-- gt3_dmonitorout_out,
      ------------------ Receive Ports - FPGA RX Interface Ports -----------------
          gt3_rxusrclk_in                 =>      gt3_rxusrclk_in,
          gt3_rxusrclk2_in                =>      gt3_rxusrclk2_in,
      ------------------ Receive Ports - FPGA RX interface Ports -----------------
          gt3_rxdata_out                  =>      gt3_rxdata_out,
      ------------------------ Receive Ports - RX AFE Ports ----------------------
          gt3_gthrxn_in                   =>       RXN_IN(3),--gt3_gthrxn_in,
      ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
          gt3_rxphmonitor_out             =>     open,-- gt3_rxphmonitor_out,
          gt3_rxphslipmonitor_out         =>    open,--  gt3_rxphslipmonitor_out,
      --------------------- Receive Ports - RX Equalizer Ports -------------------
          gt3_rxmonitorout_out            =>  open,--    gt3_rxmonitorout_out,
          gt3_rxmonitorsel_in             =>    "00",--   gt3_rxmonitorsel_in,
      --------------- Receive Ports - RX Fabric Output Control Ports -------------
          gt3_rxoutclk_out                =>      gt3_rxoutclk_out,
      ------------- Receive Ports - RX Initialization and Reset Ports ------------
          gt3_gtrxreset_in                =>      gt3_gtrxreset_in,
      ------------------------ Receive Ports -RX AFE Ports -----------------------
          gt3_gthrxp_in                   =>       RXP_IN(3),--gt3_gthrxp_in,
      -------------- Receive Ports -RX Initialization and Reset Ports ------------
          gt3_rxresetdone_out             =>      gt3_rxresetdone_out,
      --------------------- TX Initialization and Reset Ports --------------------
          gt3_gttxreset_in                =>      gt3_gttxreset_in,
          gt3_txuserrdy_in                =>      gt3_txuserrdy_in,
      ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
          gt3_txusrclk_in                 =>      gt3_txusrclk_in,
          gt3_txusrclk2_in                =>      gt3_txusrclk2_in,
      ------------------ Transmit Ports - TX Data Path interface -----------------
          gt3_txdata_in                   =>      gt3_txdata_in,
      ---------------- Transmit Ports - TX Driver and OOB signaling --------------
         gt3_gthtxn_out                  =>     TXN_OUT(3),-- gt1_gthtxn_out,
                gt3_gthtxp_out                  =>     TXP_OUT(3),-- gt1_gthtxp_out,
      ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
          gt3_txoutclk_out                =>      gt3_txoutclk_out,
          gt3_txoutclkfabric_out          =>      open,--  gt3_txoutclkfabric_out,
          gt3_txoutclkpcs_out             =>      open,--  gt3_txoutclkpcs_out,
      ------------- Transmit Ports - TX Initialization and Reset Ports -----------
          gt3_txresetdone_out             =>      gt3_txresetdone_out,
  
  
      --____________________________COMMON PORTS________________________________
       GT0_QPLLOUTCLK_IN  => '0',-- GT0_QPLLOUTCLK_IN,
       GT0_QPLLOUTREFCLK_IN => '0'--GT0_QPLLOUTREFCLK_IN 
  
  );
  




   
end RTL;


