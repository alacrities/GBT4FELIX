--Modified by Kai Chen
-- 2015/01/14
-- For FELIX: 4-chanel 4.8Gbps QPLL GTH

-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.4
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : gtwizard_qpll_4p8g_4ch.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gtwizard_qpll_4p8g_4ch (a Core Top)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************
entity gtwizard_qpll_4p8g_4ch is
generic
(
   
    STABLE_CLOCK_PERIOD                     : integer   := 24

);
port
(
    q2_clk0_refclk_in							: in   std_logic; 
   DRP_CLK_IN                            : in   std_logic;
    
    --- RX clock, for each channel
    gt0_rxusrclk_in  : in   std_logic;
    gt0_rxoutclk_out : out  std_logic;
    
    gt1_rxusrclk_in  : in   std_logic;
    gt1_rxoutclk_out : out  std_logic;
    
    gt2_rxusrclk_in  : in   std_logic;
    gt2_rxoutclk_out : out  std_logic;
    
    gt3_rxusrclk_in  : in   std_logic;
    gt3_rxoutclk_out : out  std_logic;
    
    --- TX clock, shared by all channels
    gt0_txusrclk_in    : in   std_logic;
    gt0_txoutclk_out : out  std_logic;

-----------------------------------------
---- STATUS signals
-----------------------------------------
    gt_txresetdone_out   : out  std_logic_vector(3 downto 0); 
   gt_rxresetdone_out   : out  std_logic_vector(3 downto 0);
    
    gt_txfsmresetdone_out : out  std_logic_vector(3 downto 0);
    gt_rxfsmresetdone_out : out  std_logic_vector(3 downto 0);
    
    gt_cpllfbclklost_out     : out  std_logic_vector(3 downto 0);
    gt_cplllock_out             : out  std_logic_vector(3 downto 0);
    
    gt_rxcdrlock_out         : out  std_logic_vector(3 downto 0);
    gt_qplllock_out             : out  std_logic;
---------------------------
---- CTRL signals
---------------------------
    gt_rxslide_in             : in   std_logic_vector(3 downto 0);
    gt_txuserrdy_in           : in   std_logic_vector(3 downto 0); 
    gt_rxuserrdy_in           : in   std_logic_vector(3 downto 0);
    
----------------------------------------------------------------
----------RESET SIGNALs
----------------------------------------------------------------     
    
    SOFT_RESET_IN                                   : in     std_logic; 
   GTTX_RESET_IN                           : in   std_logic_vector(3 downto 0);
   GTRX_RESET_IN                           : in   std_logic_vector(3 downto 0);
   CPLL_RESET_IN                           : in   std_logic_vector(3 downto 0);
   QPLL_RESET_IN                           : in   std_logic;
   
    SOFT_TXRST_GT      : in   std_logic_vector(3 downto 0);
      SOFT_RXRST_GT     : in   std_logic_vector(3 downto 0);
      SOFT_TXRST_ALL      : in   std_logic;
      SOFT_RXRST_ALL      : in   std_logic;

-----------------------------------------------------------
----------- Data and TX/RX Ports
-----------------------------------------------------------
    
    RX_DATA_gt0_20b : out std_logic_vector(19 downto 0);
    TX_DATA_gt0_20b : in std_logic_vector(19 downto 0);
    RX_DATA_gt1_20b : out std_logic_vector(19 downto 0);
    TX_DATA_gt1_20b : in std_logic_vector(19 downto 0);
    RX_DATA_gt2_20b : out std_logic_vector(19 downto 0);
    TX_DATA_gt2_20b : in std_logic_vector(19 downto 0);
    RX_DATA_gt3_20b : out std_logic_vector(19 downto 0);
    TX_DATA_gt3_20b : in std_logic_vector(19 downto 0);
    
   RXN_IN                                  : in   std_logic_vector(3 downto 0);
   RXP_IN                                  : in   std_logic_vector(3 downto 0);
   TXN_OUT                                 : out  std_logic_vector(3 downto 0);
   TXP_OUT                                 : out  std_logic_vector(3 downto 0)
   
   
   

);
end gtwizard_qpll_4p8g_4ch;

architecture RTL of gtwizard_qpll_4p8g_4ch is
    attribute DowngradeIPIdentifiedWarnings: string;
    attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of RTL : architecture is "gtwizard_qpll_4p8g_4ch,gtwizard_v3_4,{protocol_file=Start_from_scratch}";
    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gtwizard_qpll_4p8g_4ch,gtwizard_v3_4,{protocol_file=Start_from_scratch}";

--**************************Component Declarations*****************************

component gtwizard_qpll_4p8g_4ch_init 
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;          -- Set to 1 for simulation
 
    STABLE_CLOCK_PERIOD                     : integer   := 10;  
        -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
     SOFT_TXRST_GT      : in   std_logic_vector(3 downto 0);
            SOFT_RXRST_GT     : in   std_logic_vector(3 downto 0);
            SOFT_TXRST_ALL      : in   std_logic;
            SOFT_RXRST_ALL      : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_DRP_BUSY_OUT                        : out  std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT1_DRP_BUSY_OUT                        : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT2_DRP_BUSY_OUT                        : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT3_DRP_BUSY_OUT                        : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt0_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt0_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt0_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;

    --GT1  (X1Y5)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt1_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt1_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt1_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;

    --GT2  (X1Y6)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt2_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt2_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt2_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;

    --GT3  (X1Y7)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    --------------- Receive Ports - Comma Detection and Alignment --------------
    gt3_rxslide_in                          : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(19 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    gt3_rxphmonitor_out                     : out  std_logic_vector(4 downto 0);
    gt3_rxphslipmonitor_out                 : out  std_logic_vector(4 downto 0);
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(19 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;


    --____________________________COMMON PORTS________________________________
    GT0_QPLLLOCK_IN : in std_logic;
    GT0_QPLLREFCLKLOST_IN  : in std_logic;
    GT0_QPLLRESET_OUT  : out std_logic;
     GT0_QPLLOUTCLK_IN  : in std_logic;
     GT0_QPLLOUTREFCLK_IN : in std_logic

);
end component;

signal GT0_QPLLLOCK_I: std_logic:='0';
signal gt0_gttxreset_in : std_logic:='0';
signal gt1_gttxreset_in : std_logic:='0';
signal gt2_gttxreset_in : std_logic:='0';
signal gt3_gttxreset_in : std_logic:='0';
signal gt0_gtrxreset_in : std_logic:='0';
signal gt1_gtrxreset_in : std_logic:='0';
signal gt2_gtrxreset_in : std_logic:='0';
signal gt3_gtrxreset_in : std_logic:='0';

signal gt0_qplloutclk_i:std_logic;

 signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    
 signal gt0_drpaddr_in, gt1_drpaddr_in, gt2_drpaddr_in, gt3_drpaddr_in :  std_logic_vector(8 downto 0);   
 signal gt0_drpdi_in, gt1_drpdi_in, gt2_drpdi_in, gt3_drpdi_in :  std_logic_vector(15 downto 0);   
  signal gt0_drpdo_out, gt1_drpdo_out, gt2_drpdo_out, gt3_drpdo_out :  std_logic_vector(15 downto 0); 
  signal gt0_drpen_in, gt1_drpen_in,gt2_drpen_in,gt3_drpen_in:std_logic;
  signal gt0_drprdy_out, gt1_drprdy_out,gt2_drprdy_out,gt3_drprdy_out:std_logic;
  signal gt0_drpwe_in, gt1_drpwe_in,gt2_drpwe_in,gt3_drpwe_in:std_logic;
 signal gt1_txoutclk_out,gt2_txoutclk_out,gt3_txoutclk_out:std_logic;
 
 signal GT0_QPLLREFCLKLOST_I, GT0_QPLLRESET_I,GT0_QPLLOUTREFCLK_I:std_logic;

 
--**************************** Main Body of Code *******************************
begin

  tied_to_ground_i                             <= '0';
    tied_to_ground_vec_i                         <= x"0000000000000000";
    tied_to_vcc_i                                <= '1';
    tied_to_vcc_vec_i                            <= x"ff";


  gt_cpllfbclklost_out     <= "0000";
    gt_cplllock_out       <= "1111";
    
    gt_rxcdrlock_out        <="1111";
    gt_qplllock_out            <= GT0_QPLLLOCK_I;
   

  gt0_gttxreset_in <= GTTX_RESET_IN(0) or (not GT0_QPLLLOCK_I);
  gt1_gttxreset_in <= GTTX_RESET_IN(1) or (not GT0_QPLLLOCK_I);
  gt2_gttxreset_in <= GTTX_RESET_IN(2) or (not GT0_QPLLLOCK_I);
  gt3_gttxreset_in <= GTTX_RESET_IN(3) or (not GT0_QPLLLOCK_I);
  
  gt0_gtrxreset_in <= GTRX_RESET_IN(0) or (not GT0_QPLLLOCK_I);
  gt1_gtrxreset_in <= GTRX_RESET_IN(1) or (not GT0_QPLLLOCK_I);
  gt2_gtrxreset_in <= GTRX_RESET_IN(2) or (not GT0_QPLLLOCK_I); 
  gt3_gtrxreset_in <= GTRX_RESET_IN(3) or (not GT0_QPLLLOCK_I);



    U0 : gtwizard_qpll_4p8g_4ch_init
    generic map
(
        EXAMPLE_SIM_GTRESET_SPEEDUP   => "FALSE",
        EXAMPLE_SIMULATION            => 0,
 
        STABLE_CLOCK_PERIOD           => STABLE_CLOCK_PERIOD,
        EXAMPLE_USE_CHIPSCOPE         => 1
)
port map
(
        SYSCLK_IN                       =>      DRP_CLK_IN,
        SOFT_RESET_IN                   =>      SOFT_RESET_IN,
        
        SOFT_TXRST_GT     => SOFT_TXRST_GT,
        SOFT_RXRST_GT    => SOFT_RXRST_GT,
        SOFT_TXRST_ALL      => SOFT_TXRST_ALL,
        SOFT_RXRST_ALL     => SOFT_RXRST_ALL,
        
        DONT_RESET_ON_DATA_ERROR_IN     =>      '1',
    
    GT0_DRP_BUSY_OUT => open,
    GT0_TX_FSM_RESET_DONE_OUT => gt_txfsmresetdone_out(0),
    GT0_RX_FSM_RESET_DONE_OUT => gt_rxfsmresetdone_out(0),
    GT0_DATA_VALID_IN => '1',
    GT1_DRP_BUSY_OUT => open,
    GT1_TX_FSM_RESET_DONE_OUT => gt_txfsmresetdone_out(1),
    GT1_RX_FSM_RESET_DONE_OUT => gt_rxfsmresetdone_out(1),
    GT1_DATA_VALID_IN => '1',
    GT2_DRP_BUSY_OUT => open,
    GT2_TX_FSM_RESET_DONE_OUT => gt_txfsmresetdone_out(2),
    GT2_RX_FSM_RESET_DONE_OUT => gt_rxfsmresetdone_out(2),
    GT2_DATA_VALID_IN => '1',
    GT3_DRP_BUSY_OUT => open,
    GT3_TX_FSM_RESET_DONE_OUT => gt_txfsmresetdone_out(3),
    GT3_RX_FSM_RESET_DONE_OUT => gt_rxfsmresetdone_out(3),
    GT3_DATA_VALID_IN => '1',

    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      gt0_drpaddr_in,
        gt0_drpclk_in                   =>      DRP_CLK_IN,
        gt0_drpdi_in                    =>      gt0_drpdi_in,
        gt0_drpdo_out                   =>      gt0_drpdo_out,
        gt0_drpen_in                    =>      gt0_drpen_in,
        gt0_drprdy_out                  =>      gt0_drprdy_out,
        gt0_drpwe_in                    =>      gt0_drpwe_in,
    --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      '0',
        gt0_rxuserrdy_in                =>      gt_rxuserrdy_in(0),
    -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      open,
        gt0_eyescantrigger_in           =>      '0',
    --------------- Receive Ports - Comma Detection and Alignment --------------
        gt0_rxslide_in                  =>      gt_rxslide_in(0),
    ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt0_dmonitorout_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_in,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk_in,
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      RX_DATA_gt0_20b,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gthrxn_in                   =>      RXN_IN(0),
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt0_rxphmonitor_out             =>      open,
        gt0_rxphslipmonitor_out         =>      open,
    --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt0_rxmonitorout_out            =>      open,
        gt0_rxmonitorsel_in             =>      "00",
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_out,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_in,
    ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt0_gthrxp_in                   =>      RXP_IN(0),
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt_rxresetdone_out(0),-- gt0_rxresetdone_out,
    --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_in,
        gt0_txuserrdy_in                =>      gt_txuserrdy_in(0),
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                 =>      gt0_txusrclk_in,
        gt0_txusrclk2_in                =>      gt0_txusrclk_in,
    ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                   =>      TX_DATA_gt0_20b,
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gthtxn_out                  =>      TXN_OUT(0),
        gt0_gthtxp_out                  =>      TXP_OUT(0),
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_out,
        gt0_txoutclkfabric_out          =>      open,--gt0_txoutclkfabric_out,
        gt0_txoutclkpcs_out             =>      open,--gt0_txoutclkpcs_out,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt_txresetdone_out(0),

    --GT1  (X1Y5)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpaddr_in                  =>      gt1_drpaddr_in,
        gt1_drpclk_in                   =>      DRP_CLK_IN,
        gt1_drpdi_in                    =>      gt1_drpdi_in,
        gt1_drpdo_out                   =>      gt1_drpdo_out,
        gt1_drpen_in                    =>      gt1_drpen_in,
        gt1_drprdy_out                  =>      gt1_drprdy_out,
        gt1_drpwe_in                    =>      gt1_drpwe_in,
    --------------------- RX Initialization and Reset Ports --------------------
        gt1_eyescanreset_in             =>      '0',
        gt1_rxuserrdy_in                =>      gt_rxuserrdy_in(1),
    -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      open,
        gt1_eyescantrigger_in           =>      '0',
    --------------- Receive Ports - Comma Detection and Alignment --------------
        gt1_rxslide_in                  =>      gt_rxslide_in(1),
    ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt1_dmonitorout_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt1_rxusrclk_in,
        gt1_rxusrclk2_in                =>      gt1_rxusrclk_in,
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      RX_DATA_gt1_20b,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gthrxn_in                   =>      RXN_IN(1),
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt1_rxphmonitor_out             =>      open,
        gt1_rxphslipmonitor_out         =>      open,
    --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt1_rxmonitorout_out            =>      open,
        gt1_rxmonitorsel_in             =>      "00",
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_out,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_in,
    ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt1_gthrxp_in                   =>      RXP_IN(1),
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt_rxresetdone_out(1),
    --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_in,
        gt1_txuserrdy_in                =>      gt_txuserrdy_in(1),
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txusrclk_in                 =>      gt0_txusrclk_in,
        gt1_txusrclk2_in                =>      gt0_txusrclk_in,
    ------------------ Transmit Ports - TX Data Path interface -----------------
        gt1_txdata_in                   =>      TX_DATA_gt1_20b,
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt1_gthtxn_out                  =>      TXN_OUT(1),
        gt1_gthtxp_out                  =>      TXP_OUT(1),
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclk_out                =>      gt1_txoutclk_out,
        gt1_txoutclkfabric_out          =>      open,--gt1_txoutclkfabric_out,
        gt1_txoutclkpcs_out             =>      open,--gt1_txoutclkpcs_out,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      gt_txresetdone_out(1),

    --GT2  (X1Y6)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpaddr_in                  =>      gt2_drpaddr_in,
        gt2_drpclk_in                   =>      DRP_CLK_IN,
        gt2_drpdi_in                    =>      gt2_drpdi_in,
        gt2_drpdo_out                   =>      gt2_drpdo_out,
        gt2_drpen_in                    =>      gt2_drpen_in,
        gt2_drprdy_out                  =>      gt2_drprdy_out,
        gt2_drpwe_in                    =>      gt2_drpwe_in,
    --------------------- RX Initialization and Reset Ports --------------------
        gt2_eyescanreset_in             =>      '0',
        gt2_rxuserrdy_in                =>      gt_rxuserrdy_in(2),
    -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      open,
        gt2_eyescantrigger_in           =>      '0',
    --------------- Receive Ports - Comma Detection and Alignment --------------
        gt2_rxslide_in                  =>      gt_rxslide_in(2),
    ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt2_dmonitorout_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt2_rxusrclk_in,
        gt2_rxusrclk2_in                =>      gt2_rxusrclk_in,
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      RX_DATA_gt2_20b,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gthrxn_in                   =>      RXN_IN(2),
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt2_rxphmonitor_out             =>      open,
        gt2_rxphslipmonitor_out         =>      open,
    --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt2_rxmonitorout_out            =>      open,
        gt2_rxmonitorsel_in             =>      "00",
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_out,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_in,
    ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt2_gthrxp_in                   =>      RXP_IN(2),
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt_rxresetdone_out(2),
    --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_in,
        gt2_txuserrdy_in                =>      gt_txuserrdy_in(2),
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txusrclk_in                 =>      gt0_txusrclk_in,
        gt2_txusrclk2_in                =>      gt0_txusrclk_in,
    ------------------ Transmit Ports - TX Data Path interface -----------------
        gt2_txdata_in                   =>      TX_DATA_gt2_20b,
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt2_gthtxn_out                  =>      TXN_OUT(2),
        gt2_gthtxp_out                  =>      TXP_OUT(2),
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclk_out                =>      gt2_txoutclk_out,
        gt2_txoutclkfabric_out          =>      open,--gt2_txoutclkfabric_out,
        gt2_txoutclkpcs_out             =>      open,--gt2_txoutclkpcs_out,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      gt_txresetdone_out(2),

    --GT3  (X1Y7)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpaddr_in                  =>      gt3_drpaddr_in,
        gt3_drpclk_in                   =>      DRP_CLK_IN,
        gt3_drpdi_in                    =>      gt3_drpdi_in,
        gt3_drpdo_out                   =>      gt3_drpdo_out,
        gt3_drpen_in                    =>      gt3_drpen_in,
        gt3_drprdy_out                  =>      gt3_drprdy_out,
        gt3_drpwe_in                    =>      gt3_drpwe_in,
    --------------------- RX Initialization and Reset Ports --------------------
        gt3_eyescanreset_in             =>      '0',
        gt3_rxuserrdy_in                =>      gt_rxuserrdy_in(3),
    -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      open,
        gt3_eyescantrigger_in           =>      '0',
    --------------- Receive Ports - Comma Detection and Alignment --------------
        gt3_rxslide_in                  =>      gt_rxslide_in(3),
    ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt3_dmonitorout_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt3_rxusrclk_in,
        gt3_rxusrclk2_in                =>      gt3_rxusrclk_in,
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      RX_DATA_gt3_20b,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gthrxn_in                   =>      RXN_IN(3),
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        gt3_rxphmonitor_out             =>      open,
        gt3_rxphslipmonitor_out         =>      open,
    --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt3_rxmonitorout_out            =>      open,
        gt3_rxmonitorsel_in             =>      "00",
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_out,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_in,
    ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt3_gthrxp_in                   =>      RXP_IN(3),
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt_rxresetdone_out(3),
    --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_in,
        gt3_txuserrdy_in                =>      gt_txuserrdy_in(3),
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txusrclk_in                 =>      gt0_txusrclk_in,
        gt3_txusrclk2_in                =>      gt0_txusrclk_in,
    ------------------ Transmit Ports - TX Data Path interface -----------------
        gt3_txdata_in                   =>      TX_DATA_gt3_20b,
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt3_gthtxn_out                  =>      TXN_OUT(3),
        gt3_gthtxp_out                  =>      TXP_OUT(3),
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclk_out                =>      gt3_txoutclk_out,
        gt3_txoutclkfabric_out          =>      open,--gt3_txoutclkfabric_out,
        gt3_txoutclkpcs_out             =>      open,--gt3_txoutclkpcs_out,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      gt_txresetdone_out(3),


    --____________________________COMMON PORTS________________________________
    GT0_QPLLLOCK_IN => GT0_QPLLLOCK_I, 
    GT0_QPLLREFCLKLOST_IN => GT0_QPLLREFCLKLOST_I, 
    GT0_QPLLRESET_OUT => GT0_QPLLRESET_I, 
     GT0_QPLLOUTCLK_IN  => GT0_QPLLOUTCLK_I,
     GT0_QPLLOUTREFCLK_IN => GT0_QPLLOUTREFCLK_I 

);

    gthe2_common_0_i : GTHE2_COMMON
    generic map
    (
            -- Simulation attributes
            SIM_RESET_SPEEDUP    => ("FALSE"),
            SIM_QPLLREFCLK_SEL   => ("001"),
            SIM_VERSION          => ("2.0"),


       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000040000001050"),
        COMMON_CFG                              =>     (x"0000001C"),
        QPLL_CFG                                =>     (x"04801C7"),
        QPLL_CLKOUT_CFG                         =>     ("1111"),
        QPLL_COARSE_FREQ_OVRD                   =>     ("010000"),
        QPLL_COARSE_FREQ_OVRD_EN                =>     ('0'),
        QPLL_CP                                 =>     ("0000011111"),
        QPLL_CP_MONITOR_EN                      =>     ('0'),
        QPLL_DMONITOR_SEL                       =>     ('0'),
        QPLL_FBDIV                              =>     ("0010000000"),--(QPLL_FBDIV_IN),
        QPLL_FBDIV_MONITOR_EN                   =>     ('0'),
        QPLL_FBDIV_RATIO                        =>      ('1'),--(QPLL_FBDIV_RATIO),
        QPLL_INIT_CFG                           =>     (x"000006"),
        QPLL_LOCK_CFG                           =>     (x"05E8"),
        QPLL_LPF                                =>     ("1111"),
        QPLL_REFCLK_DIV                         =>     (1),
        RSVD_ATTR0                              =>     (x"0000"),
        RSVD_ATTR1                              =>     (x"0000"),
        QPLL_RP_COMP                            =>     ('0'),
        QPLL_VTRL_RESET                         =>     ("00"),
        RCAL_CFG                                =>     ("00")

        
    )
    port map
    (
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GTGREFCLK                       =>      tied_to_ground_i,
        GTNORTHREFCLK0                  =>      tied_to_ground_i,
        GTNORTHREFCLK1                  =>      tied_to_ground_i,
        GTREFCLK0                       =>      q2_clk0_refclk_in,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTSOUTHREFCLK0                  =>      tied_to_ground_i,
        GTSOUTHREFCLK1                  =>      tied_to_ground_i,
        ------------------------- Common Block -  QPLL Ports -----------------------
        QPLLDMONITOR                    =>      open,
        ----------------------- Common Block - Clocking Ports ----------------------
        QPLLOUTCLK                      =>      gt0_qplloutclk_i,
        QPLLOUTREFCLK                   =>      gt0_qplloutrefclk_i,
        REFCLKOUTMONITOR                =>      open,
        ------------------------- Common Block - QPLL Ports ------------------------
        BGRCALOVRDENB                   =>      tied_to_vcc_i,
        PMARSVDOUT                      =>      open,
        QPLLFBCLKLOST                   =>      open,
        QPLLLOCK                        =>      GT0_QPLLLOCK_I,
        QPLLLOCKDETCLK                  =>      DRP_CLK_IN,
        QPLLLOCKEN                      =>      tied_to_vcc_i,
        QPLLOUTRESET                    =>      tied_to_ground_i,
        QPLLPD                          =>      tied_to_ground_i,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_I,
        QPLLREFCLKSEL                   =>      "001",
        QPLLRESET                       =>      GT0_QPLLRESET_i or QPLL_RESET_IN,
        QPLLRSVD1                       =>      "0000000000000000",
        QPLLRSVD2                       =>      "11111",
        --------------------------------- QPLL Ports -------------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i

    );


 
end RTL;    
 
